module timer1hz_tb ();

  reg clk_100MHz, reset;
  wire clk_1Hz;


endmodule
